module sectioner

pub struct Config {

}